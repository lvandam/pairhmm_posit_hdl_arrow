../../../../pairhmm_posit_hdl/pairhmm/Sources/afu/rtl/pe.vhd