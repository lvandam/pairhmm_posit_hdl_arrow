../../../../pairhmm_posit_hdl/pairhmm/Sources/afu/rtl/pairhmm.vhd